magic
tech sky130A
magscale 1 2
timestamp 1636340147
<< obsli1 >>
rect 1104 1105 244323 244273
<< obsm1 >>
rect 658 960 244335 244304
<< metal2 >>
rect 1030 245869 1086 246669
rect 3146 245869 3202 246669
rect 5262 245869 5318 246669
rect 7378 245869 7434 246669
rect 9586 245869 9642 246669
rect 11702 245869 11758 246669
rect 13818 245869 13874 246669
rect 16026 245869 16082 246669
rect 18142 245869 18198 246669
rect 20258 245869 20314 246669
rect 22466 245869 22522 246669
rect 24582 245869 24638 246669
rect 26698 245869 26754 246669
rect 28906 245869 28962 246669
rect 31022 245869 31078 246669
rect 33138 245869 33194 246669
rect 35346 245869 35402 246669
rect 37462 245869 37518 246669
rect 39578 245869 39634 246669
rect 41786 245869 41842 246669
rect 43902 245869 43958 246669
rect 46018 245869 46074 246669
rect 48134 245869 48190 246669
rect 50342 245869 50398 246669
rect 52458 245869 52514 246669
rect 54574 245869 54630 246669
rect 56782 245869 56838 246669
rect 58898 245869 58954 246669
rect 61014 245869 61070 246669
rect 63222 245869 63278 246669
rect 65338 245869 65394 246669
rect 67454 245869 67510 246669
rect 69662 245869 69718 246669
rect 71778 245869 71834 246669
rect 73894 245869 73950 246669
rect 76102 245869 76158 246669
rect 78218 245869 78274 246669
rect 80334 245869 80390 246669
rect 82542 245869 82598 246669
rect 84658 245869 84714 246669
rect 86774 245869 86830 246669
rect 88890 245869 88946 246669
rect 91098 245869 91154 246669
rect 93214 245869 93270 246669
rect 95330 245869 95386 246669
rect 97538 245869 97594 246669
rect 99654 245869 99710 246669
rect 101770 245869 101826 246669
rect 103978 245869 104034 246669
rect 106094 245869 106150 246669
rect 108210 245869 108266 246669
rect 110418 245869 110474 246669
rect 112534 245869 112590 246669
rect 114650 245869 114706 246669
rect 116858 245869 116914 246669
rect 118974 245869 119030 246669
rect 121090 245869 121146 246669
rect 123298 245869 123354 246669
rect 125414 245869 125470 246669
rect 127530 245869 127586 246669
rect 129646 245869 129702 246669
rect 131854 245869 131910 246669
rect 133970 245869 134026 246669
rect 136086 245869 136142 246669
rect 138294 245869 138350 246669
rect 140410 245869 140466 246669
rect 142526 245869 142582 246669
rect 144734 245869 144790 246669
rect 146850 245869 146906 246669
rect 148966 245869 149022 246669
rect 151174 245869 151230 246669
rect 153290 245869 153346 246669
rect 155406 245869 155462 246669
rect 157614 245869 157670 246669
rect 159730 245869 159786 246669
rect 161846 245869 161902 246669
rect 164054 245869 164110 246669
rect 166170 245869 166226 246669
rect 168286 245869 168342 246669
rect 170402 245869 170458 246669
rect 172610 245869 172666 246669
rect 174726 245869 174782 246669
rect 176842 245869 176898 246669
rect 179050 245869 179106 246669
rect 181166 245869 181222 246669
rect 183282 245869 183338 246669
rect 185490 245869 185546 246669
rect 187606 245869 187662 246669
rect 189722 245869 189778 246669
rect 191930 245869 191986 246669
rect 194046 245869 194102 246669
rect 196162 245869 196218 246669
rect 198370 245869 198426 246669
rect 200486 245869 200542 246669
rect 202602 245869 202658 246669
rect 204810 245869 204866 246669
rect 206926 245869 206982 246669
rect 209042 245869 209098 246669
rect 211158 245869 211214 246669
rect 213366 245869 213422 246669
rect 215482 245869 215538 246669
rect 217598 245869 217654 246669
rect 219806 245869 219862 246669
rect 221922 245869 221978 246669
rect 224038 245869 224094 246669
rect 226246 245869 226302 246669
rect 228362 245869 228418 246669
rect 230478 245869 230534 246669
rect 232686 245869 232742 246669
rect 234802 245869 234858 246669
rect 236918 245869 236974 246669
rect 239126 245869 239182 246669
rect 241242 245869 241298 246669
rect 243358 245869 243414 246669
rect 202 0 258 800
rect 662 0 718 800
rect 1122 0 1178 800
rect 1674 0 1730 800
rect 2134 0 2190 800
rect 2594 0 2650 800
rect 3146 0 3202 800
rect 3606 0 3662 800
rect 4158 0 4214 800
rect 4618 0 4674 800
rect 5078 0 5134 800
rect 5630 0 5686 800
rect 6090 0 6146 800
rect 6642 0 6698 800
rect 7102 0 7158 800
rect 7562 0 7618 800
rect 8114 0 8170 800
rect 8574 0 8630 800
rect 9126 0 9182 800
rect 9586 0 9642 800
rect 10046 0 10102 800
rect 10598 0 10654 800
rect 11058 0 11114 800
rect 11610 0 11666 800
rect 12070 0 12126 800
rect 12530 0 12586 800
rect 13082 0 13138 800
rect 13542 0 13598 800
rect 14002 0 14058 800
rect 14554 0 14610 800
rect 15014 0 15070 800
rect 15566 0 15622 800
rect 16026 0 16082 800
rect 16486 0 16542 800
rect 17038 0 17094 800
rect 17498 0 17554 800
rect 18050 0 18106 800
rect 18510 0 18566 800
rect 18970 0 19026 800
rect 19522 0 19578 800
rect 19982 0 20038 800
rect 20534 0 20590 800
rect 20994 0 21050 800
rect 21454 0 21510 800
rect 22006 0 22062 800
rect 22466 0 22522 800
rect 23018 0 23074 800
rect 23478 0 23534 800
rect 23938 0 23994 800
rect 24490 0 24546 800
rect 24950 0 25006 800
rect 25410 0 25466 800
rect 25962 0 26018 800
rect 26422 0 26478 800
rect 26974 0 27030 800
rect 27434 0 27490 800
rect 27894 0 27950 800
rect 28446 0 28502 800
rect 28906 0 28962 800
rect 29458 0 29514 800
rect 29918 0 29974 800
rect 30378 0 30434 800
rect 30930 0 30986 800
rect 31390 0 31446 800
rect 31942 0 31998 800
rect 32402 0 32458 800
rect 32862 0 32918 800
rect 33414 0 33470 800
rect 33874 0 33930 800
rect 34426 0 34482 800
rect 34886 0 34942 800
rect 35346 0 35402 800
rect 35898 0 35954 800
rect 36358 0 36414 800
rect 36818 0 36874 800
rect 37370 0 37426 800
rect 37830 0 37886 800
rect 38382 0 38438 800
rect 38842 0 38898 800
rect 39302 0 39358 800
rect 39854 0 39910 800
rect 40314 0 40370 800
rect 40866 0 40922 800
rect 41326 0 41382 800
rect 41786 0 41842 800
rect 42338 0 42394 800
rect 42798 0 42854 800
rect 43350 0 43406 800
rect 43810 0 43866 800
rect 44270 0 44326 800
rect 44822 0 44878 800
rect 45282 0 45338 800
rect 45834 0 45890 800
rect 46294 0 46350 800
rect 46754 0 46810 800
rect 47306 0 47362 800
rect 47766 0 47822 800
rect 48226 0 48282 800
rect 48778 0 48834 800
rect 49238 0 49294 800
rect 49790 0 49846 800
rect 50250 0 50306 800
rect 50710 0 50766 800
rect 51262 0 51318 800
rect 51722 0 51778 800
rect 52274 0 52330 800
rect 52734 0 52790 800
rect 53194 0 53250 800
rect 53746 0 53802 800
rect 54206 0 54262 800
rect 54758 0 54814 800
rect 55218 0 55274 800
rect 55678 0 55734 800
rect 56230 0 56286 800
rect 56690 0 56746 800
rect 57242 0 57298 800
rect 57702 0 57758 800
rect 58162 0 58218 800
rect 58714 0 58770 800
rect 59174 0 59230 800
rect 59634 0 59690 800
rect 60186 0 60242 800
rect 60646 0 60702 800
rect 61198 0 61254 800
rect 61658 0 61714 800
rect 62118 0 62174 800
rect 62670 0 62726 800
rect 63130 0 63186 800
rect 63682 0 63738 800
rect 64142 0 64198 800
rect 64602 0 64658 800
rect 65154 0 65210 800
rect 65614 0 65670 800
rect 66166 0 66222 800
rect 66626 0 66682 800
rect 67086 0 67142 800
rect 67638 0 67694 800
rect 68098 0 68154 800
rect 68650 0 68706 800
rect 69110 0 69166 800
rect 69570 0 69626 800
rect 70122 0 70178 800
rect 70582 0 70638 800
rect 71042 0 71098 800
rect 71594 0 71650 800
rect 72054 0 72110 800
rect 72606 0 72662 800
rect 73066 0 73122 800
rect 73526 0 73582 800
rect 74078 0 74134 800
rect 74538 0 74594 800
rect 75090 0 75146 800
rect 75550 0 75606 800
rect 76010 0 76066 800
rect 76562 0 76618 800
rect 77022 0 77078 800
rect 77574 0 77630 800
rect 78034 0 78090 800
rect 78494 0 78550 800
rect 79046 0 79102 800
rect 79506 0 79562 800
rect 80058 0 80114 800
rect 80518 0 80574 800
rect 80978 0 81034 800
rect 81530 0 81586 800
rect 81990 0 82046 800
rect 82450 0 82506 800
rect 83002 0 83058 800
rect 83462 0 83518 800
rect 84014 0 84070 800
rect 84474 0 84530 800
rect 84934 0 84990 800
rect 85486 0 85542 800
rect 85946 0 86002 800
rect 86498 0 86554 800
rect 86958 0 87014 800
rect 87418 0 87474 800
rect 87970 0 88026 800
rect 88430 0 88486 800
rect 88982 0 89038 800
rect 89442 0 89498 800
rect 89902 0 89958 800
rect 90454 0 90510 800
rect 90914 0 90970 800
rect 91466 0 91522 800
rect 91926 0 91982 800
rect 92386 0 92442 800
rect 92938 0 92994 800
rect 93398 0 93454 800
rect 93858 0 93914 800
rect 94410 0 94466 800
rect 94870 0 94926 800
rect 95422 0 95478 800
rect 95882 0 95938 800
rect 96342 0 96398 800
rect 96894 0 96950 800
rect 97354 0 97410 800
rect 97906 0 97962 800
rect 98366 0 98422 800
rect 98826 0 98882 800
rect 99378 0 99434 800
rect 99838 0 99894 800
rect 100390 0 100446 800
rect 100850 0 100906 800
rect 101310 0 101366 800
rect 101862 0 101918 800
rect 102322 0 102378 800
rect 102874 0 102930 800
rect 103334 0 103390 800
rect 103794 0 103850 800
rect 104346 0 104402 800
rect 104806 0 104862 800
rect 105266 0 105322 800
rect 105818 0 105874 800
rect 106278 0 106334 800
rect 106830 0 106886 800
rect 107290 0 107346 800
rect 107750 0 107806 800
rect 108302 0 108358 800
rect 108762 0 108818 800
rect 109314 0 109370 800
rect 109774 0 109830 800
rect 110234 0 110290 800
rect 110786 0 110842 800
rect 111246 0 111302 800
rect 111798 0 111854 800
rect 112258 0 112314 800
rect 112718 0 112774 800
rect 113270 0 113326 800
rect 113730 0 113786 800
rect 114282 0 114338 800
rect 114742 0 114798 800
rect 115202 0 115258 800
rect 115754 0 115810 800
rect 116214 0 116270 800
rect 116674 0 116730 800
rect 117226 0 117282 800
rect 117686 0 117742 800
rect 118238 0 118294 800
rect 118698 0 118754 800
rect 119158 0 119214 800
rect 119710 0 119766 800
rect 120170 0 120226 800
rect 120722 0 120778 800
rect 121182 0 121238 800
rect 121642 0 121698 800
rect 122194 0 122250 800
rect 122654 0 122710 800
rect 123206 0 123262 800
rect 123666 0 123722 800
rect 124126 0 124182 800
rect 124678 0 124734 800
rect 125138 0 125194 800
rect 125690 0 125746 800
rect 126150 0 126206 800
rect 126610 0 126666 800
rect 127162 0 127218 800
rect 127622 0 127678 800
rect 128174 0 128230 800
rect 128634 0 128690 800
rect 129094 0 129150 800
rect 129646 0 129702 800
rect 130106 0 130162 800
rect 130566 0 130622 800
rect 131118 0 131174 800
rect 131578 0 131634 800
rect 132130 0 132186 800
rect 132590 0 132646 800
rect 133050 0 133106 800
rect 133602 0 133658 800
rect 134062 0 134118 800
rect 134614 0 134670 800
rect 135074 0 135130 800
rect 135534 0 135590 800
rect 136086 0 136142 800
rect 136546 0 136602 800
rect 137098 0 137154 800
rect 137558 0 137614 800
rect 138018 0 138074 800
rect 138570 0 138626 800
rect 139030 0 139086 800
rect 139582 0 139638 800
rect 140042 0 140098 800
rect 140502 0 140558 800
rect 141054 0 141110 800
rect 141514 0 141570 800
rect 141974 0 142030 800
rect 142526 0 142582 800
rect 142986 0 143042 800
rect 143538 0 143594 800
rect 143998 0 144054 800
rect 144458 0 144514 800
rect 145010 0 145066 800
rect 145470 0 145526 800
rect 146022 0 146078 800
rect 146482 0 146538 800
rect 146942 0 146998 800
rect 147494 0 147550 800
rect 147954 0 148010 800
rect 148506 0 148562 800
rect 148966 0 149022 800
rect 149426 0 149482 800
rect 149978 0 150034 800
rect 150438 0 150494 800
rect 150990 0 151046 800
rect 151450 0 151506 800
rect 151910 0 151966 800
rect 152462 0 152518 800
rect 152922 0 152978 800
rect 153382 0 153438 800
rect 153934 0 153990 800
rect 154394 0 154450 800
rect 154946 0 155002 800
rect 155406 0 155462 800
rect 155866 0 155922 800
rect 156418 0 156474 800
rect 156878 0 156934 800
rect 157430 0 157486 800
rect 157890 0 157946 800
rect 158350 0 158406 800
rect 158902 0 158958 800
rect 159362 0 159418 800
rect 159914 0 159970 800
rect 160374 0 160430 800
rect 160834 0 160890 800
rect 161386 0 161442 800
rect 161846 0 161902 800
rect 162398 0 162454 800
rect 162858 0 162914 800
rect 163318 0 163374 800
rect 163870 0 163926 800
rect 164330 0 164386 800
rect 164790 0 164846 800
rect 165342 0 165398 800
rect 165802 0 165858 800
rect 166354 0 166410 800
rect 166814 0 166870 800
rect 167274 0 167330 800
rect 167826 0 167882 800
rect 168286 0 168342 800
rect 168838 0 168894 800
rect 169298 0 169354 800
rect 169758 0 169814 800
rect 170310 0 170366 800
rect 170770 0 170826 800
rect 171322 0 171378 800
rect 171782 0 171838 800
rect 172242 0 172298 800
rect 172794 0 172850 800
rect 173254 0 173310 800
rect 173806 0 173862 800
rect 174266 0 174322 800
rect 174726 0 174782 800
rect 175278 0 175334 800
rect 175738 0 175794 800
rect 176198 0 176254 800
rect 176750 0 176806 800
rect 177210 0 177266 800
rect 177762 0 177818 800
rect 178222 0 178278 800
rect 178682 0 178738 800
rect 179234 0 179290 800
rect 179694 0 179750 800
rect 180246 0 180302 800
rect 180706 0 180762 800
rect 181166 0 181222 800
rect 181718 0 181774 800
rect 182178 0 182234 800
rect 182730 0 182786 800
rect 183190 0 183246 800
rect 183650 0 183706 800
rect 184202 0 184258 800
rect 184662 0 184718 800
rect 185214 0 185270 800
rect 185674 0 185730 800
rect 186134 0 186190 800
rect 186686 0 186742 800
rect 187146 0 187202 800
rect 187606 0 187662 800
rect 188158 0 188214 800
rect 188618 0 188674 800
rect 189170 0 189226 800
rect 189630 0 189686 800
rect 190090 0 190146 800
rect 190642 0 190698 800
rect 191102 0 191158 800
rect 191654 0 191710 800
rect 192114 0 192170 800
rect 192574 0 192630 800
rect 193126 0 193182 800
rect 193586 0 193642 800
rect 194138 0 194194 800
rect 194598 0 194654 800
rect 195058 0 195114 800
rect 195610 0 195666 800
rect 196070 0 196126 800
rect 196622 0 196678 800
rect 197082 0 197138 800
rect 197542 0 197598 800
rect 198094 0 198150 800
rect 198554 0 198610 800
rect 199014 0 199070 800
rect 199566 0 199622 800
rect 200026 0 200082 800
rect 200578 0 200634 800
rect 201038 0 201094 800
rect 201498 0 201554 800
rect 202050 0 202106 800
rect 202510 0 202566 800
rect 203062 0 203118 800
rect 203522 0 203578 800
rect 203982 0 204038 800
rect 204534 0 204590 800
rect 204994 0 205050 800
rect 205546 0 205602 800
rect 206006 0 206062 800
rect 206466 0 206522 800
rect 207018 0 207074 800
rect 207478 0 207534 800
rect 208030 0 208086 800
rect 208490 0 208546 800
rect 208950 0 209006 800
rect 209502 0 209558 800
rect 209962 0 210018 800
rect 210422 0 210478 800
rect 210974 0 211030 800
rect 211434 0 211490 800
rect 211986 0 212042 800
rect 212446 0 212502 800
rect 212906 0 212962 800
rect 213458 0 213514 800
rect 213918 0 213974 800
rect 214470 0 214526 800
rect 214930 0 214986 800
rect 215390 0 215446 800
rect 215942 0 215998 800
rect 216402 0 216458 800
rect 216954 0 217010 800
rect 217414 0 217470 800
rect 217874 0 217930 800
rect 218426 0 218482 800
rect 218886 0 218942 800
rect 219438 0 219494 800
rect 219898 0 219954 800
rect 220358 0 220414 800
rect 220910 0 220966 800
rect 221370 0 221426 800
rect 221830 0 221886 800
rect 222382 0 222438 800
rect 222842 0 222898 800
rect 223394 0 223450 800
rect 223854 0 223910 800
rect 224314 0 224370 800
rect 224866 0 224922 800
rect 225326 0 225382 800
rect 225878 0 225934 800
rect 226338 0 226394 800
rect 226798 0 226854 800
rect 227350 0 227406 800
rect 227810 0 227866 800
rect 228362 0 228418 800
rect 228822 0 228878 800
rect 229282 0 229338 800
rect 229834 0 229890 800
rect 230294 0 230350 800
rect 230846 0 230902 800
rect 231306 0 231362 800
rect 231766 0 231822 800
rect 232318 0 232374 800
rect 232778 0 232834 800
rect 233238 0 233294 800
rect 233790 0 233846 800
rect 234250 0 234306 800
rect 234802 0 234858 800
rect 235262 0 235318 800
rect 235722 0 235778 800
rect 236274 0 236330 800
rect 236734 0 236790 800
rect 237286 0 237342 800
rect 237746 0 237802 800
rect 238206 0 238262 800
rect 238758 0 238814 800
rect 239218 0 239274 800
rect 239770 0 239826 800
rect 240230 0 240286 800
rect 240690 0 240746 800
rect 241242 0 241298 800
rect 241702 0 241758 800
rect 242254 0 242310 800
rect 242714 0 242770 800
rect 243174 0 243230 800
rect 243726 0 243782 800
rect 244186 0 244242 800
<< obsm2 >>
rect 202 245813 974 245869
rect 1142 245813 3090 245869
rect 3258 245813 5206 245869
rect 5374 245813 7322 245869
rect 7490 245813 9530 245869
rect 9698 245813 11646 245869
rect 11814 245813 13762 245869
rect 13930 245813 15970 245869
rect 16138 245813 18086 245869
rect 18254 245813 20202 245869
rect 20370 245813 22410 245869
rect 22578 245813 24526 245869
rect 24694 245813 26642 245869
rect 26810 245813 28850 245869
rect 29018 245813 30966 245869
rect 31134 245813 33082 245869
rect 33250 245813 35290 245869
rect 35458 245813 37406 245869
rect 37574 245813 39522 245869
rect 39690 245813 41730 245869
rect 41898 245813 43846 245869
rect 44014 245813 45962 245869
rect 46130 245813 48078 245869
rect 48246 245813 50286 245869
rect 50454 245813 52402 245869
rect 52570 245813 54518 245869
rect 54686 245813 56726 245869
rect 56894 245813 58842 245869
rect 59010 245813 60958 245869
rect 61126 245813 63166 245869
rect 63334 245813 65282 245869
rect 65450 245813 67398 245869
rect 67566 245813 69606 245869
rect 69774 245813 71722 245869
rect 71890 245813 73838 245869
rect 74006 245813 76046 245869
rect 76214 245813 78162 245869
rect 78330 245813 80278 245869
rect 80446 245813 82486 245869
rect 82654 245813 84602 245869
rect 84770 245813 86718 245869
rect 86886 245813 88834 245869
rect 89002 245813 91042 245869
rect 91210 245813 93158 245869
rect 93326 245813 95274 245869
rect 95442 245813 97482 245869
rect 97650 245813 99598 245869
rect 99766 245813 101714 245869
rect 101882 245813 103922 245869
rect 104090 245813 106038 245869
rect 106206 245813 108154 245869
rect 108322 245813 110362 245869
rect 110530 245813 112478 245869
rect 112646 245813 114594 245869
rect 114762 245813 116802 245869
rect 116970 245813 118918 245869
rect 119086 245813 121034 245869
rect 121202 245813 123242 245869
rect 123410 245813 125358 245869
rect 125526 245813 127474 245869
rect 127642 245813 129590 245869
rect 129758 245813 131798 245869
rect 131966 245813 133914 245869
rect 134082 245813 136030 245869
rect 136198 245813 138238 245869
rect 138406 245813 140354 245869
rect 140522 245813 142470 245869
rect 142638 245813 144678 245869
rect 144846 245813 146794 245869
rect 146962 245813 148910 245869
rect 149078 245813 151118 245869
rect 151286 245813 153234 245869
rect 153402 245813 155350 245869
rect 155518 245813 157558 245869
rect 157726 245813 159674 245869
rect 159842 245813 161790 245869
rect 161958 245813 163998 245869
rect 164166 245813 166114 245869
rect 166282 245813 168230 245869
rect 168398 245813 170346 245869
rect 170514 245813 172554 245869
rect 172722 245813 174670 245869
rect 174838 245813 176786 245869
rect 176954 245813 178994 245869
rect 179162 245813 181110 245869
rect 181278 245813 183226 245869
rect 183394 245813 185434 245869
rect 185602 245813 187550 245869
rect 187718 245813 189666 245869
rect 189834 245813 191874 245869
rect 192042 245813 193990 245869
rect 194158 245813 196106 245869
rect 196274 245813 198314 245869
rect 198482 245813 200430 245869
rect 200598 245813 202546 245869
rect 202714 245813 204754 245869
rect 204922 245813 206870 245869
rect 207038 245813 208986 245869
rect 209154 245813 211102 245869
rect 211270 245813 213310 245869
rect 213478 245813 215426 245869
rect 215594 245813 217542 245869
rect 217710 245813 219750 245869
rect 219918 245813 221866 245869
rect 222034 245813 223982 245869
rect 224150 245813 226190 245869
rect 226358 245813 228306 245869
rect 228474 245813 230422 245869
rect 230590 245813 232630 245869
rect 232798 245813 234746 245869
rect 234914 245813 236862 245869
rect 237030 245813 239070 245869
rect 239238 245813 241186 245869
rect 241354 245813 243302 245869
rect 243470 245813 244240 245869
rect 202 856 244240 245813
rect 314 734 606 856
rect 774 734 1066 856
rect 1234 734 1618 856
rect 1786 734 2078 856
rect 2246 734 2538 856
rect 2706 734 3090 856
rect 3258 734 3550 856
rect 3718 734 4102 856
rect 4270 734 4562 856
rect 4730 734 5022 856
rect 5190 734 5574 856
rect 5742 734 6034 856
rect 6202 734 6586 856
rect 6754 734 7046 856
rect 7214 734 7506 856
rect 7674 734 8058 856
rect 8226 734 8518 856
rect 8686 734 9070 856
rect 9238 734 9530 856
rect 9698 734 9990 856
rect 10158 734 10542 856
rect 10710 734 11002 856
rect 11170 734 11554 856
rect 11722 734 12014 856
rect 12182 734 12474 856
rect 12642 734 13026 856
rect 13194 734 13486 856
rect 13654 734 13946 856
rect 14114 734 14498 856
rect 14666 734 14958 856
rect 15126 734 15510 856
rect 15678 734 15970 856
rect 16138 734 16430 856
rect 16598 734 16982 856
rect 17150 734 17442 856
rect 17610 734 17994 856
rect 18162 734 18454 856
rect 18622 734 18914 856
rect 19082 734 19466 856
rect 19634 734 19926 856
rect 20094 734 20478 856
rect 20646 734 20938 856
rect 21106 734 21398 856
rect 21566 734 21950 856
rect 22118 734 22410 856
rect 22578 734 22962 856
rect 23130 734 23422 856
rect 23590 734 23882 856
rect 24050 734 24434 856
rect 24602 734 24894 856
rect 25062 734 25354 856
rect 25522 734 25906 856
rect 26074 734 26366 856
rect 26534 734 26918 856
rect 27086 734 27378 856
rect 27546 734 27838 856
rect 28006 734 28390 856
rect 28558 734 28850 856
rect 29018 734 29402 856
rect 29570 734 29862 856
rect 30030 734 30322 856
rect 30490 734 30874 856
rect 31042 734 31334 856
rect 31502 734 31886 856
rect 32054 734 32346 856
rect 32514 734 32806 856
rect 32974 734 33358 856
rect 33526 734 33818 856
rect 33986 734 34370 856
rect 34538 734 34830 856
rect 34998 734 35290 856
rect 35458 734 35842 856
rect 36010 734 36302 856
rect 36470 734 36762 856
rect 36930 734 37314 856
rect 37482 734 37774 856
rect 37942 734 38326 856
rect 38494 734 38786 856
rect 38954 734 39246 856
rect 39414 734 39798 856
rect 39966 734 40258 856
rect 40426 734 40810 856
rect 40978 734 41270 856
rect 41438 734 41730 856
rect 41898 734 42282 856
rect 42450 734 42742 856
rect 42910 734 43294 856
rect 43462 734 43754 856
rect 43922 734 44214 856
rect 44382 734 44766 856
rect 44934 734 45226 856
rect 45394 734 45778 856
rect 45946 734 46238 856
rect 46406 734 46698 856
rect 46866 734 47250 856
rect 47418 734 47710 856
rect 47878 734 48170 856
rect 48338 734 48722 856
rect 48890 734 49182 856
rect 49350 734 49734 856
rect 49902 734 50194 856
rect 50362 734 50654 856
rect 50822 734 51206 856
rect 51374 734 51666 856
rect 51834 734 52218 856
rect 52386 734 52678 856
rect 52846 734 53138 856
rect 53306 734 53690 856
rect 53858 734 54150 856
rect 54318 734 54702 856
rect 54870 734 55162 856
rect 55330 734 55622 856
rect 55790 734 56174 856
rect 56342 734 56634 856
rect 56802 734 57186 856
rect 57354 734 57646 856
rect 57814 734 58106 856
rect 58274 734 58658 856
rect 58826 734 59118 856
rect 59286 734 59578 856
rect 59746 734 60130 856
rect 60298 734 60590 856
rect 60758 734 61142 856
rect 61310 734 61602 856
rect 61770 734 62062 856
rect 62230 734 62614 856
rect 62782 734 63074 856
rect 63242 734 63626 856
rect 63794 734 64086 856
rect 64254 734 64546 856
rect 64714 734 65098 856
rect 65266 734 65558 856
rect 65726 734 66110 856
rect 66278 734 66570 856
rect 66738 734 67030 856
rect 67198 734 67582 856
rect 67750 734 68042 856
rect 68210 734 68594 856
rect 68762 734 69054 856
rect 69222 734 69514 856
rect 69682 734 70066 856
rect 70234 734 70526 856
rect 70694 734 70986 856
rect 71154 734 71538 856
rect 71706 734 71998 856
rect 72166 734 72550 856
rect 72718 734 73010 856
rect 73178 734 73470 856
rect 73638 734 74022 856
rect 74190 734 74482 856
rect 74650 734 75034 856
rect 75202 734 75494 856
rect 75662 734 75954 856
rect 76122 734 76506 856
rect 76674 734 76966 856
rect 77134 734 77518 856
rect 77686 734 77978 856
rect 78146 734 78438 856
rect 78606 734 78990 856
rect 79158 734 79450 856
rect 79618 734 80002 856
rect 80170 734 80462 856
rect 80630 734 80922 856
rect 81090 734 81474 856
rect 81642 734 81934 856
rect 82102 734 82394 856
rect 82562 734 82946 856
rect 83114 734 83406 856
rect 83574 734 83958 856
rect 84126 734 84418 856
rect 84586 734 84878 856
rect 85046 734 85430 856
rect 85598 734 85890 856
rect 86058 734 86442 856
rect 86610 734 86902 856
rect 87070 734 87362 856
rect 87530 734 87914 856
rect 88082 734 88374 856
rect 88542 734 88926 856
rect 89094 734 89386 856
rect 89554 734 89846 856
rect 90014 734 90398 856
rect 90566 734 90858 856
rect 91026 734 91410 856
rect 91578 734 91870 856
rect 92038 734 92330 856
rect 92498 734 92882 856
rect 93050 734 93342 856
rect 93510 734 93802 856
rect 93970 734 94354 856
rect 94522 734 94814 856
rect 94982 734 95366 856
rect 95534 734 95826 856
rect 95994 734 96286 856
rect 96454 734 96838 856
rect 97006 734 97298 856
rect 97466 734 97850 856
rect 98018 734 98310 856
rect 98478 734 98770 856
rect 98938 734 99322 856
rect 99490 734 99782 856
rect 99950 734 100334 856
rect 100502 734 100794 856
rect 100962 734 101254 856
rect 101422 734 101806 856
rect 101974 734 102266 856
rect 102434 734 102818 856
rect 102986 734 103278 856
rect 103446 734 103738 856
rect 103906 734 104290 856
rect 104458 734 104750 856
rect 104918 734 105210 856
rect 105378 734 105762 856
rect 105930 734 106222 856
rect 106390 734 106774 856
rect 106942 734 107234 856
rect 107402 734 107694 856
rect 107862 734 108246 856
rect 108414 734 108706 856
rect 108874 734 109258 856
rect 109426 734 109718 856
rect 109886 734 110178 856
rect 110346 734 110730 856
rect 110898 734 111190 856
rect 111358 734 111742 856
rect 111910 734 112202 856
rect 112370 734 112662 856
rect 112830 734 113214 856
rect 113382 734 113674 856
rect 113842 734 114226 856
rect 114394 734 114686 856
rect 114854 734 115146 856
rect 115314 734 115698 856
rect 115866 734 116158 856
rect 116326 734 116618 856
rect 116786 734 117170 856
rect 117338 734 117630 856
rect 117798 734 118182 856
rect 118350 734 118642 856
rect 118810 734 119102 856
rect 119270 734 119654 856
rect 119822 734 120114 856
rect 120282 734 120666 856
rect 120834 734 121126 856
rect 121294 734 121586 856
rect 121754 734 122138 856
rect 122306 734 122598 856
rect 122766 734 123150 856
rect 123318 734 123610 856
rect 123778 734 124070 856
rect 124238 734 124622 856
rect 124790 734 125082 856
rect 125250 734 125634 856
rect 125802 734 126094 856
rect 126262 734 126554 856
rect 126722 734 127106 856
rect 127274 734 127566 856
rect 127734 734 128118 856
rect 128286 734 128578 856
rect 128746 734 129038 856
rect 129206 734 129590 856
rect 129758 734 130050 856
rect 130218 734 130510 856
rect 130678 734 131062 856
rect 131230 734 131522 856
rect 131690 734 132074 856
rect 132242 734 132534 856
rect 132702 734 132994 856
rect 133162 734 133546 856
rect 133714 734 134006 856
rect 134174 734 134558 856
rect 134726 734 135018 856
rect 135186 734 135478 856
rect 135646 734 136030 856
rect 136198 734 136490 856
rect 136658 734 137042 856
rect 137210 734 137502 856
rect 137670 734 137962 856
rect 138130 734 138514 856
rect 138682 734 138974 856
rect 139142 734 139526 856
rect 139694 734 139986 856
rect 140154 734 140446 856
rect 140614 734 140998 856
rect 141166 734 141458 856
rect 141626 734 141918 856
rect 142086 734 142470 856
rect 142638 734 142930 856
rect 143098 734 143482 856
rect 143650 734 143942 856
rect 144110 734 144402 856
rect 144570 734 144954 856
rect 145122 734 145414 856
rect 145582 734 145966 856
rect 146134 734 146426 856
rect 146594 734 146886 856
rect 147054 734 147438 856
rect 147606 734 147898 856
rect 148066 734 148450 856
rect 148618 734 148910 856
rect 149078 734 149370 856
rect 149538 734 149922 856
rect 150090 734 150382 856
rect 150550 734 150934 856
rect 151102 734 151394 856
rect 151562 734 151854 856
rect 152022 734 152406 856
rect 152574 734 152866 856
rect 153034 734 153326 856
rect 153494 734 153878 856
rect 154046 734 154338 856
rect 154506 734 154890 856
rect 155058 734 155350 856
rect 155518 734 155810 856
rect 155978 734 156362 856
rect 156530 734 156822 856
rect 156990 734 157374 856
rect 157542 734 157834 856
rect 158002 734 158294 856
rect 158462 734 158846 856
rect 159014 734 159306 856
rect 159474 734 159858 856
rect 160026 734 160318 856
rect 160486 734 160778 856
rect 160946 734 161330 856
rect 161498 734 161790 856
rect 161958 734 162342 856
rect 162510 734 162802 856
rect 162970 734 163262 856
rect 163430 734 163814 856
rect 163982 734 164274 856
rect 164442 734 164734 856
rect 164902 734 165286 856
rect 165454 734 165746 856
rect 165914 734 166298 856
rect 166466 734 166758 856
rect 166926 734 167218 856
rect 167386 734 167770 856
rect 167938 734 168230 856
rect 168398 734 168782 856
rect 168950 734 169242 856
rect 169410 734 169702 856
rect 169870 734 170254 856
rect 170422 734 170714 856
rect 170882 734 171266 856
rect 171434 734 171726 856
rect 171894 734 172186 856
rect 172354 734 172738 856
rect 172906 734 173198 856
rect 173366 734 173750 856
rect 173918 734 174210 856
rect 174378 734 174670 856
rect 174838 734 175222 856
rect 175390 734 175682 856
rect 175850 734 176142 856
rect 176310 734 176694 856
rect 176862 734 177154 856
rect 177322 734 177706 856
rect 177874 734 178166 856
rect 178334 734 178626 856
rect 178794 734 179178 856
rect 179346 734 179638 856
rect 179806 734 180190 856
rect 180358 734 180650 856
rect 180818 734 181110 856
rect 181278 734 181662 856
rect 181830 734 182122 856
rect 182290 734 182674 856
rect 182842 734 183134 856
rect 183302 734 183594 856
rect 183762 734 184146 856
rect 184314 734 184606 856
rect 184774 734 185158 856
rect 185326 734 185618 856
rect 185786 734 186078 856
rect 186246 734 186630 856
rect 186798 734 187090 856
rect 187258 734 187550 856
rect 187718 734 188102 856
rect 188270 734 188562 856
rect 188730 734 189114 856
rect 189282 734 189574 856
rect 189742 734 190034 856
rect 190202 734 190586 856
rect 190754 734 191046 856
rect 191214 734 191598 856
rect 191766 734 192058 856
rect 192226 734 192518 856
rect 192686 734 193070 856
rect 193238 734 193530 856
rect 193698 734 194082 856
rect 194250 734 194542 856
rect 194710 734 195002 856
rect 195170 734 195554 856
rect 195722 734 196014 856
rect 196182 734 196566 856
rect 196734 734 197026 856
rect 197194 734 197486 856
rect 197654 734 198038 856
rect 198206 734 198498 856
rect 198666 734 198958 856
rect 199126 734 199510 856
rect 199678 734 199970 856
rect 200138 734 200522 856
rect 200690 734 200982 856
rect 201150 734 201442 856
rect 201610 734 201994 856
rect 202162 734 202454 856
rect 202622 734 203006 856
rect 203174 734 203466 856
rect 203634 734 203926 856
rect 204094 734 204478 856
rect 204646 734 204938 856
rect 205106 734 205490 856
rect 205658 734 205950 856
rect 206118 734 206410 856
rect 206578 734 206962 856
rect 207130 734 207422 856
rect 207590 734 207974 856
rect 208142 734 208434 856
rect 208602 734 208894 856
rect 209062 734 209446 856
rect 209614 734 209906 856
rect 210074 734 210366 856
rect 210534 734 210918 856
rect 211086 734 211378 856
rect 211546 734 211930 856
rect 212098 734 212390 856
rect 212558 734 212850 856
rect 213018 734 213402 856
rect 213570 734 213862 856
rect 214030 734 214414 856
rect 214582 734 214874 856
rect 215042 734 215334 856
rect 215502 734 215886 856
rect 216054 734 216346 856
rect 216514 734 216898 856
rect 217066 734 217358 856
rect 217526 734 217818 856
rect 217986 734 218370 856
rect 218538 734 218830 856
rect 218998 734 219382 856
rect 219550 734 219842 856
rect 220010 734 220302 856
rect 220470 734 220854 856
rect 221022 734 221314 856
rect 221482 734 221774 856
rect 221942 734 222326 856
rect 222494 734 222786 856
rect 222954 734 223338 856
rect 223506 734 223798 856
rect 223966 734 224258 856
rect 224426 734 224810 856
rect 224978 734 225270 856
rect 225438 734 225822 856
rect 225990 734 226282 856
rect 226450 734 226742 856
rect 226910 734 227294 856
rect 227462 734 227754 856
rect 227922 734 228306 856
rect 228474 734 228766 856
rect 228934 734 229226 856
rect 229394 734 229778 856
rect 229946 734 230238 856
rect 230406 734 230790 856
rect 230958 734 231250 856
rect 231418 734 231710 856
rect 231878 734 232262 856
rect 232430 734 232722 856
rect 232890 734 233182 856
rect 233350 734 233734 856
rect 233902 734 234194 856
rect 234362 734 234746 856
rect 234914 734 235206 856
rect 235374 734 235666 856
rect 235834 734 236218 856
rect 236386 734 236678 856
rect 236846 734 237230 856
rect 237398 734 237690 856
rect 237858 734 238150 856
rect 238318 734 238702 856
rect 238870 734 239162 856
rect 239330 734 239714 856
rect 239882 734 240174 856
rect 240342 734 240634 856
rect 240802 734 241186 856
rect 241354 734 241646 856
rect 241814 734 242198 856
rect 242366 734 242658 856
rect 242826 734 243118 856
rect 243286 734 243670 856
rect 243838 734 244130 856
<< obsm3 >>
rect 197 1667 243235 244289
<< metal4 >>
rect 4208 2128 4528 244304
rect 19568 2128 19888 244304
rect 34928 2128 35248 244304
rect 50288 2128 50608 244304
rect 65648 2128 65968 244304
rect 81008 2128 81328 244304
rect 96368 2128 96688 244304
rect 111728 2128 112048 244304
rect 127088 2128 127408 244304
rect 142448 2128 142768 244304
rect 157808 2128 158128 244304
rect 173168 2128 173488 244304
rect 188528 2128 188848 244304
rect 203888 2128 204208 244304
rect 219248 2128 219568 244304
rect 234608 2128 234928 244304
<< obsm4 >>
rect 2635 2048 4128 240141
rect 4608 2048 19488 240141
rect 19968 2048 34848 240141
rect 35328 2048 50208 240141
rect 50688 2048 65568 240141
rect 66048 2048 80928 240141
rect 81408 2048 96288 240141
rect 96768 2048 111648 240141
rect 112128 2048 127008 240141
rect 127488 2048 142368 240141
rect 142848 2048 157728 240141
rect 158208 2048 173088 240141
rect 173568 2048 188448 240141
rect 188928 2048 203808 240141
rect 204288 2048 219168 240141
rect 219648 2048 234528 240141
rect 235008 2048 239693 240141
rect 2635 1939 239693 2048
<< labels >>
rlabel metal2 s 1030 245869 1086 246669 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 65338 245869 65394 246669 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 71778 245869 71834 246669 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 78218 245869 78274 246669 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 84658 245869 84714 246669 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 91098 245869 91154 246669 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 97538 245869 97594 246669 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 103978 245869 104034 246669 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 110418 245869 110474 246669 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 116858 245869 116914 246669 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 123298 245869 123354 246669 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 7378 245869 7434 246669 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 129646 245869 129702 246669 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 136086 245869 136142 246669 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 142526 245869 142582 246669 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 148966 245869 149022 246669 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 155406 245869 155462 246669 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 161846 245869 161902 246669 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 168286 245869 168342 246669 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 174726 245869 174782 246669 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 181166 245869 181222 246669 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 187606 245869 187662 246669 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 13818 245869 13874 246669 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 194046 245869 194102 246669 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 200486 245869 200542 246669 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 206926 245869 206982 246669 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 213366 245869 213422 246669 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 219806 245869 219862 246669 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 226246 245869 226302 246669 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 232686 245869 232742 246669 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 239126 245869 239182 246669 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 20258 245869 20314 246669 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 26698 245869 26754 246669 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 33138 245869 33194 246669 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 39578 245869 39634 246669 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 46018 245869 46074 246669 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 52458 245869 52514 246669 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 58898 245869 58954 246669 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3146 245869 3202 246669 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 67454 245869 67510 246669 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 73894 245869 73950 246669 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 80334 245869 80390 246669 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 86774 245869 86830 246669 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 93214 245869 93270 246669 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 99654 245869 99710 246669 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 106094 245869 106150 246669 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 112534 245869 112590 246669 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 118974 245869 119030 246669 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 125414 245869 125470 246669 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 9586 245869 9642 246669 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 131854 245869 131910 246669 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 138294 245869 138350 246669 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 144734 245869 144790 246669 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 151174 245869 151230 246669 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 157614 245869 157670 246669 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 164054 245869 164110 246669 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 170402 245869 170458 246669 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 176842 245869 176898 246669 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 183282 245869 183338 246669 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 189722 245869 189778 246669 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 16026 245869 16082 246669 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 196162 245869 196218 246669 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 202602 245869 202658 246669 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 209042 245869 209098 246669 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 215482 245869 215538 246669 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 221922 245869 221978 246669 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 228362 245869 228418 246669 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 234802 245869 234858 246669 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 241242 245869 241298 246669 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 22466 245869 22522 246669 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 28906 245869 28962 246669 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 35346 245869 35402 246669 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 41786 245869 41842 246669 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 48134 245869 48190 246669 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 54574 245869 54630 246669 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 61014 245869 61070 246669 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 5262 245869 5318 246669 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 69662 245869 69718 246669 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 76102 245869 76158 246669 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 82542 245869 82598 246669 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 88890 245869 88946 246669 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 95330 245869 95386 246669 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 101770 245869 101826 246669 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 108210 245869 108266 246669 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 114650 245869 114706 246669 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 121090 245869 121146 246669 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 127530 245869 127586 246669 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 11702 245869 11758 246669 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 133970 245869 134026 246669 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 140410 245869 140466 246669 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 146850 245869 146906 246669 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 153290 245869 153346 246669 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 159730 245869 159786 246669 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 166170 245869 166226 246669 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 172610 245869 172666 246669 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 179050 245869 179106 246669 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 185490 245869 185546 246669 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 191930 245869 191986 246669 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 18142 245869 18198 246669 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 198370 245869 198426 246669 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 204810 245869 204866 246669 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 211158 245869 211214 246669 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 217598 245869 217654 246669 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 224038 245869 224094 246669 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 230478 245869 230534 246669 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 236918 245869 236974 246669 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 243358 245869 243414 246669 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 24582 245869 24638 246669 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 31022 245869 31078 246669 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 37462 245869 37518 246669 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 43902 245869 43958 246669 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 50342 245869 50398 246669 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 56782 245869 56838 246669 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 63222 245869 63278 246669 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 243174 0 243230 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 243726 0 243782 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 244186 0 244242 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 52734 0 52790 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 201498 0 201554 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 203062 0 203118 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 204534 0 204590 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 206006 0 206062 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 207478 0 207534 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 208950 0 209006 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 210422 0 210478 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 211986 0 212042 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 213458 0 213514 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 214930 0 214986 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 216402 0 216458 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 217874 0 217930 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 219438 0 219494 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 220910 0 220966 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 222382 0 222438 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 223854 0 223910 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 225326 0 225382 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 226798 0 226854 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 228362 0 228418 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 229834 0 229890 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 231306 0 231362 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 232778 0 232834 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 234250 0 234306 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 235722 0 235778 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 237286 0 237342 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 238758 0 238814 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 240230 0 240286 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 241702 0 241758 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 76562 0 76618 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 78034 0 78090 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 79506 0 79562 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 97354 0 97410 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 101862 0 101918 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 103334 0 103390 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 107750 0 107806 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 109314 0 109370 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 110786 0 110842 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 112258 0 112314 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 113730 0 113786 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 115202 0 115258 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 116674 0 116730 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 118238 0 118294 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 119710 0 119766 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 121182 0 121238 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 124126 0 124182 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 127162 0 127218 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 128634 0 128690 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 133050 0 133106 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 134614 0 134670 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 136086 0 136142 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 137558 0 137614 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 139030 0 139086 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 140502 0 140558 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 141974 0 142030 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 143538 0 143594 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 145010 0 145066 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 146482 0 146538 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 147954 0 148010 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 149426 0 149482 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 150990 0 151046 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 152462 0 152518 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 153934 0 153990 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 155406 0 155462 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 156878 0 156934 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 158350 0 158406 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 159914 0 159970 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 161386 0 161442 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 162858 0 162914 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 164330 0 164386 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 165802 0 165858 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 167274 0 167330 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 168838 0 168894 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 170310 0 170366 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 171782 0 171838 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 173254 0 173310 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 174726 0 174782 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 176198 0 176254 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 177762 0 177818 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 179234 0 179290 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 180706 0 180762 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 182178 0 182234 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 183650 0 183706 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 185214 0 185270 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 186686 0 186742 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 188158 0 188214 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 189630 0 189686 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 191102 0 191158 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 192574 0 192630 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 194138 0 194194 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 195610 0 195666 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 197082 0 197138 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 198554 0 198610 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 200026 0 200082 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 202050 0 202106 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 203522 0 203578 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 204994 0 205050 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 206466 0 206522 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 208030 0 208086 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 209502 0 209558 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 210974 0 211030 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 212446 0 212502 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 213918 0 213974 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 215390 0 215446 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 68098 0 68154 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 216954 0 217010 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 218426 0 218482 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 219898 0 219954 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 221370 0 221426 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 222842 0 222898 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 224314 0 224370 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 225878 0 225934 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 227350 0 227406 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 228822 0 228878 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 230294 0 230350 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 231766 0 231822 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 233238 0 233294 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 234802 0 234858 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 236274 0 236330 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 237746 0 237802 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 239218 0 239274 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 240690 0 240746 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 242254 0 242310 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 71042 0 71098 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 72606 0 72662 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 75550 0 75606 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 77022 0 77078 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 78494 0 78550 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 80058 0 80114 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 81530 0 81586 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 83002 0 83058 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 84474 0 84530 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 85946 0 86002 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 87418 0 87474 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 88982 0 89038 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 90454 0 90510 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 91926 0 91982 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 94870 0 94926 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 96342 0 96398 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 97906 0 97962 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 99378 0 99434 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 100850 0 100906 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 102322 0 102378 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 103794 0 103850 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 105266 0 105322 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 108302 0 108358 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 109774 0 109830 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 111246 0 111302 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 57702 0 57758 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 114282 0 114338 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 115754 0 115810 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 117226 0 117282 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 118698 0 118754 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 120170 0 120226 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 121642 0 121698 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 123206 0 123262 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 124678 0 124734 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 126150 0 126206 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 59174 0 59230 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 127622 0 127678 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 129094 0 129150 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 130566 0 130622 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 132130 0 132186 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 133602 0 133658 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 135074 0 135130 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 136546 0 136602 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 138018 0 138074 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 139582 0 139638 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 141054 0 141110 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 60646 0 60702 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 142526 0 142582 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 143998 0 144054 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 145470 0 145526 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 146942 0 146998 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 148506 0 148562 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 149978 0 150034 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 151450 0 151506 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 152922 0 152978 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 154394 0 154450 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 155866 0 155922 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 62118 0 62174 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 157430 0 157486 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 158902 0 158958 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 160374 0 160430 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 161846 0 161902 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 163318 0 163374 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 164790 0 164846 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 166354 0 166410 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 167826 0 167882 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 169298 0 169354 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 170770 0 170826 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 63682 0 63738 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 172242 0 172298 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 173806 0 173862 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 175278 0 175334 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 176750 0 176806 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 178222 0 178278 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 179694 0 179750 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 181166 0 181222 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 182730 0 182786 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 184202 0 184258 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 185674 0 185730 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 65154 0 65210 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 187146 0 187202 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 188618 0 188674 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 190090 0 190146 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 191654 0 191710 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 193126 0 193182 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 194598 0 194654 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 196070 0 196126 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 197542 0 197598 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 199014 0 199070 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 200578 0 200634 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 66626 0 66682 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 53746 0 53802 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 202510 0 202566 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 203982 0 204038 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 205546 0 205602 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 207018 0 207074 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 208490 0 208546 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 209962 0 210018 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 211434 0 211490 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 212906 0 212962 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 214470 0 214526 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 215942 0 215998 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 217414 0 217470 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 218886 0 218942 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 220358 0 220414 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 221830 0 221886 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 223394 0 223450 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 224866 0 224922 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 226338 0 226394 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 227810 0 227866 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 229282 0 229338 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 230846 0 230902 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 232318 0 232374 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 233790 0 233846 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 235262 0 235318 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 236734 0 236790 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 238206 0 238262 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 239770 0 239826 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 241242 0 241298 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 242714 0 242770 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 89442 0 89498 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 101310 0 101366 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 108762 0 108818 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 110234 0 110290 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 111798 0 111854 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 113270 0 113326 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 116214 0 116270 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 117686 0 117742 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 122194 0 122250 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 125138 0 125194 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 126610 0 126666 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 128174 0 128230 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 129646 0 129702 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 131118 0 131174 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 132590 0 132646 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 134062 0 134118 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 137098 0 137154 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 138570 0 138626 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 140042 0 140098 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 141514 0 141570 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 142986 0 143042 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 144458 0 144514 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 146022 0 146078 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 147494 0 147550 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 148966 0 149022 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 150438 0 150494 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 151910 0 151966 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 153382 0 153438 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 154946 0 155002 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 156418 0 156474 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 157890 0 157946 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 159362 0 159418 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 160834 0 160890 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 162398 0 162454 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 163870 0 163926 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 165342 0 165398 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 166814 0 166870 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 168286 0 168342 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 169758 0 169814 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 171322 0 171378 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 172794 0 172850 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 174266 0 174322 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 175738 0 175794 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 177210 0 177266 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 178682 0 178738 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 180246 0 180302 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 181718 0 181774 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 183190 0 183246 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 184662 0 184718 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 186134 0 186190 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 187606 0 187662 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 189170 0 189226 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 190642 0 190698 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 192114 0 192170 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 193586 0 193642 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 195058 0 195114 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 196622 0 196678 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 198094 0 198150 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 199566 0 199622 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 201038 0 201094 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 67086 0 67142 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 244304 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 244304 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 244304 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 244304 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 244304 6 vccd1
port 502 nsew power input
rlabel metal4 s 157808 2128 158128 244304 6 vccd1
port 502 nsew power input
rlabel metal4 s 188528 2128 188848 244304 6 vccd1
port 502 nsew power input
rlabel metal4 s 219248 2128 219568 244304 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 244304 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 244304 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 244304 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 244304 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 244304 6 vssd1
port 503 nsew ground input
rlabel metal4 s 173168 2128 173488 244304 6 vssd1
port 503 nsew ground input
rlabel metal4 s 203888 2128 204208 244304 6 vssd1
port 503 nsew ground input
rlabel metal4 s 234608 2128 234928 244304 6 vssd1
port 503 nsew ground input
rlabel metal2 s 202 0 258 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 662 0 718 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 3146 0 3202 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 28446 0 28502 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 29918 0 29974 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 6090 0 6146 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 35898 0 35954 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 38842 0 38898 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 40314 0 40370 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 41786 0 41842 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 43350 0 43406 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 44822 0 44878 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 46294 0 46350 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 47766 0 47822 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 49238 0 49294 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 8114 0 8170 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 50710 0 50766 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 52274 0 52330 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 10046 0 10102 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 12070 0 12126 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 15014 0 15070 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 4618 0 4674 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 244525 246669
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 133889676
string GDS_START 1257614
<< end >>

